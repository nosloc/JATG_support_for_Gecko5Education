`timescale 1ns/1ps

module tb_clock_synchronizer;

    // Testbench signals
    reg clk_in;
    reg clk_out;
    reg[9:0] to_sync;
    reg n_reset;
    wire[9:0] sync_out;

    // Instantiate the DUT (Device Under Test)
    clock_synchronizer #(10) uut (
        .clk_in(clk_in),
        .clk_out(clk_out),
        .to_sync(to_sync),
        .sync_out(sync_out),
        .n_reset(n_reset)
    );

    // Clock generation for clk_in
    initial begin
        clk_in = 0;
        forever #5 clk_in = ~clk_in; // 10ns period
    end

    // Clock generation for clk_out
    initial begin
        clk_out = 0;
        forever #7 clk_out = ~clk_out; // 14ns period
    end

    // Test stimulus
    initial begin
        // Initialize inputs
        to_sync = 0; // Set to_sync high
        n_reset = 0;
        #10 n_reset = 1; // Release reset after 10ns


        #10 to_sync = 10'h3FF;

        // Finish simulation
        #100 $finish;
    end

    // Monitor signals
    initial begin
         $dumpfile("test_clock_sync.vcd");
        $dumpvars(0, tb_clock_synchronizer);
    end

endmodule